code 
<!DOCTYPE sv>
	<sv>
	<head>
	<title>Page Title</title>
	</head>
	<body>
	 <h1>This is a Heading</h1>
         <p>this is a system.</p>
	  
	 </body>
	 </sv>

